module NOTgate(z,a);
  input a;
  output z;
  not#1(z,a);
endmodule